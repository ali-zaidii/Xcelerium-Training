package alu_pkg;

    typedef enum logic [2:0] {
        ADD,
        SUB,
        AND_OP,
        OR_OP,
        XOR_OP,
        SHIFT_LEFT,
        SHIFT_RIGHT
    } alu_op_t;

endpackage

